LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODE_COMPARATOR IS 
	PORT(
		DATA1  : in STD_LOGIC_VECTOR(31 downto 0);
		DATA2  : in STD_LOGIC_VECTOR(31 DOWNTO 0);
		DATAOUT: OUT STD_LOGIC
	);
END DECODE_COMPARATOR;

ARCHITECTURE BEHAVIOUR OF DECODE_COMPARATOR IS 

BEGIN 

	PROCESS (DATA1,DATA2)
		BEGIN
			IF DATA1 = DATA2 THEN
				DATAOUT <= '1';
			ELSE 
				DATAOUT <= '0';
        END IF;
    END PROCESS;
	
END BEHAVIOUR;